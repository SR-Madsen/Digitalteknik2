library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SinusKurve is
    Port ( Xakse : in STD_LOGIC_VECTOR (9 downto 0);
           xfunc : in STD_LOGIC;
           Yakse : out STD_LOGIC_VECTOR (8 downto 0));
end SinusKurve;

architecture Behavioral of SinusKurve is
    signal Sin: integer := 0;
begin   
    process( Xakse)
		variable vAdr: integer;
		variable vSin: integer;
    begin	
        if xfunc='1' then
            vAdr := conv_integer( Xakse(7 downto 0));
            if vAdr>127 then
                vAdr := 255-vAdr;
            end if;
        else
           vAdr := conv_integer( Xakse);
        end if;
		
        case vAdr is
            when 0  => vSin := 127;
            when 1  => vSin := 129;
            when 2  => vSin := 130;
            when 3  => vSin := 132;
            when 4  => vSin := 133;
            when 5  => vSin := 135;
            when 6  => vSin := 136;
            when 7  => vSin := 138;
            when 8  => vSin := 139;
            when 9  => vSin :=141;
            when 10 => vSin :=143;
            when 11 => vSin :=144;
            when 12 => vSin :=146;
            when 13 => vSin :=147;
            when 14 => vSin :=149;
            when 15 => vSin :=150;
            when 16 => vSin :=152;
            when 17 => vSin :=153;
            when 18 => vSin :=155;
            when 19 => vSin :=156;
            when 20 => vSin :=158;
            when 21 => vSin :=159;
            when 22 => vSin :=161;
            when 23 => vSin :=162;
            when 24 => vSin :=164;
            when 25 => vSin :=165;
            when 26 => vSin :=167;
            when 27 => vSin :=168;
            when 28 => vSin :=170;
            when 29 => vSin :=171;
            when 30 => vSin :=173;
            when 31 => vSin :=174;
            when 32 => vSin :=176;
            when 33 => vSin :=177;
            when 34 => vSin :=178;
            when 35 => vSin :=180;
            when 36 => vSin :=181;
            when 37 => vSin :=183;
            when 38 => vSin :=184;
            when 39 => vSin :=185;
            when 40 => vSin :=187;
            when 41 => vSin :=188;
            when 42 =>  vSin :=190;
            when 43 =>  vSin :=191;
            when 44 =>  vSin :=192;		
            when 45 =>  vSin :=194; 
            when 46 =>  vSin :=195;
            when 47 =>  vSin :=196;
            when 48 =>  vSin :=198;
            when 49 =>  vSin :=199;
            when 50 =>  vSin :=200;
            when 51 =>  vSin :=201;
            when 52 =>  vSin :=203;
            when 53 =>  vSin :=204;
            when 54 =>  vSin :=205;
            when 55 =>  vSin :=206;
            when 56 =>  vSin :=208;
            when 57 =>  vSin :=209;
            when 58 =>  vSin :=210;
            when 59 =>  vSin :=211;
            when 60 =>  vSin :=212;
            when 61 =>  vSin :=213;
            when 62 =>  vSin :=215;
            when 63 =>  vSin :=216;
            when 64 =>  vSin :=217;
            when 65 =>  vSin :=218;
            when 66 =>  vSin :=219;
            when 67 =>  vSin :=220;
            when 68 =>  vSin :=221;
            when 69 =>  vSin :=222;
            when 70 =>  vSin :=223;
            when 71 =>  vSin :=224;
            when 72 =>  vSin :=225;
            when 73 =>  vSin :=226;
            when 74 =>  vSin :=227;
            when 75 =>  vSin :=228;
            when 76 =>  vSin :=229;
            when 77 =>  vSin :=230;
            when 78 =>  vSin :=231;
            when 79 =>  vSin :=232;
            when 80 =>  vSin :=233;
            when 81 =>  vSin :=233;
            when 82 =>  vSin :=234;
            when 83 =>  vSin :=235;
            when 84 =>  vSin :=236;
            when 85 =>  vSin :=237;
            when 86 =>  vSin :=238;
            when 87 =>  vSin :=238;
            when 88 =>  vSin :=239;
            when 89 =>  vSin :=240;
            when 90 =>  vSin :=240;
            when 91 =>  vSin :=241;
            when 92 =>  vSin :=242;
            when 93 =>  vSin :=242;
            when 94 =>  vSin :=243;
            when 95 =>  vSin :=244;
            when 96 =>  vSin :=244;
            when 97 =>  vSin :=245;
            when 98 =>  vSin :=245;
            when 99 =>  vSin :=246;
            when 100 => vSin :=247;
            when 101 => vSin :=247;
            when 102 => vSin :=248;
            when 103 => vSin :=248;
            when 104 => vSin :=249;
            when 105 => vSin :=249;
            when 106 => vSin :=249;
            when 107 => vSin :=250;
            when 108 => vSin :=250;
            when 109 => vSin :=251;
            when 110 => vSin :=251;
            when 111 => vSin :=251;
            when 112 => vSin :=252;
            when 113 => vSin :=252;
            when 114 => vSin :=252;
            when 115 => vSin :=252;
            when 116 => vSin :=253;
            when 117 => vSin :=253;
            when 118 => vSin :=253;
            when 119 => vSin :=253;
            when 120 => vSin :=253;
            when 121 => vSin :=254;
            when 122 => vSin :=254;
            when 123 => vSin :=254;
            when 124 => vSin :=254;
            when 125 => vSin :=254;
            when 126 => vSin :=254;
            when 127 => vSin :=254;
            when others => vSin  := 255;
		end case;
	    
	    Yakse <= conv_std_logic_vector( vSin,9);	
    end process;
end Behavioral;
